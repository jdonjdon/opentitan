// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class chip_sw_pwm_pulses_vseq extends chip_sw_base_vseq;
  `uvm_object_utils(chip_sw_pwm_pulses_vseq)

  `uvm_object_new
 
  virtual task body();
    super.body();
    
    `uvm_info(`gfn, "Not implemented", UVM_LOW)  
  endtask // body
   
endclass // chip_sw_pwm_pulses_vseq
